library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

package parametros is

		constant n : natural:=8;
		constant m : natural:=4;

end package parametros;

package body parametros is

end;
